library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
 
package util_pkg is
 
	subtype sl is std_logic;
	subtype slv is std_logic_vector;
	type aslv is array(integer range <>) of slv;

  type state_t is (s_idle, s_detect_preamble, s_read_dst_mac, s_read_src_mac, s_read_len, s_read_data, s_get_crc);
  type ll_state_t is (s_idle, s_send_preamble, s_send_dst_mac, s_send_src_mac, s_send_len, s_send_data, s_send_crc);
  type ROM is array (natural range <>) of std_logic_vector(7 downto 0);
	function log2c(n : integer) return integer;

 
  constant etherTraff: ROM(0 to 8191) := (
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AB", x"EC", x"FF", x"44", x"47", x"45",
  x"D8", x"56", x"A4", x"89", x"EF", x"13", x"49", x"00", x"5F", x"96", x"CF", x"1A", x"A9", x"0B", x"62", x"01", x"94", x"38", x"D0", x"DA", x"51", x"68", x"4A", x"22", x"BC",
  x"8F", x"CB", x"C5", x"93", x"A5", x"01", x"E1", x"FC", x"24", x"A1", x"6D", x"00", x"E9", x"0B", x"D8", x"63", x"97", x"F5", x"74", x"D7", x"83", x"9A", x"46", x"DF", x"BB",
  x"97", x"87", x"BA", x"AC", x"C0", x"F8", x"2A", x"B4", x"09", x"49", x"13", x"AF", x"2A", x"0B", x"A7", x"93", x"FF", x"4A", x"CD", x"78", x"E4", x"98", x"98", x"89", x"09",
  x"7D", x"0D", x"D2", x"3A", x"11", x"18", x"D2", x"B3", x"1D", x"7C", x"40", x"5C", x"6E", x"7F", x"A6", x"C6", x"E2", x"DD", x"94", x"0A", x"C7", x"3E", x"D4", x"A5", x"96",
  x"96", x"3E", x"F1", x"AA", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"AA", x"AA", x"AA", x"AA", x"AA",
  x"AA", x"AA", x"AB", x"3A", x"77", x"37", x"2F", x"20", x"D0", x"15", x"AD", x"4F", x"33", x"EF", x"1F", x"00", x"54", x"C0", x"EE", x"39", x"EA", x"79", x"C4", x"5B", x"C6",
  x"11", x"2F", x"11", x"05", x"18", x"95", x"8A", x"15", x"F8", x"D2", x"A6", x"6D", x"51", x"C5", x"C9", x"7F", x"9E", x"52", x"54", x"52", x"F9", x"27", x"6D", x"92", x"70",
  x"09", x"E1", x"EA", x"32", x"0A", x"1A", x"9E", x"B8", x"5C", x"D1", x"68", x"79", x"09", x"54", x"D5", x"CA", x"06", x"44", x"2A", x"6A", x"AA", x"81", x"4F", x"B5", x"BC",
  x"55", x"B4", x"C6", x"E5", x"0E", x"6D", x"97", x"11", x"07", x"22", x"4D", x"68", x"84", x"90", x"36", x"2F", x"7E", x"51", x"E1", x"38", x"F7", x"E0", x"45", x"49", x"CA",
  x"55", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AB",
  x"E2", x"AA", x"64", x"03", x"BC", x"12", x"2B", x"FB", x"2F", x"6E", x"55", x"E0", x"00", x"32", x"CC", x"A7", x"91", x"79", x"38", x"96", x"10", x"3C", x"FA", x"8F", x"A5",
  x"7D", x"C9", x"9A", x"2E", x"55", x"0E", x"1F", x"2E", x"C4", x"EF", x"1E", x"BD", x"F8", x"A6", x"5F", x"95", x"3D", x"58", x"76", x"15", x"9B", x"C0", x"49", x"26", x"C5",
  x"85", x"D4", x"96", x"35", x"23", x"1E", x"C0", x"29", x"6C", x"C0", x"1C", x"CA", x"6C", x"25", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AB", x"DA", x"EE", x"FF", x"49", x"2D", x"94", x"0B", x"94", x"A1", x"02", x"CF", x"A2",
  x"00", x"35", x"B1", x"B1", x"BA", x"5C", x"4A", x"1B", x"1E", x"40", x"AC", x"0C", x"8E", x"56", x"C8", x"AB", x"57", x"C3", x"56", x"F4", x"D5", x"2B", x"F4", x"6D", x"67",
  x"BD", x"8D", x"B3", x"D9", x"A5", x"08", x"0A", x"93", x"DC", x"7A", x"99", x"DD", x"3D", x"45", x"11", x"E1", x"7D", x"85", x"32", x"E2", x"96", x"75", x"F9", x"76", x"5E",
  x"87", x"5B", x"63", x"87", x"CE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"AA", x"AA", x"AA", x"AA",
  x"AA", x"AA", x"AA", x"AB", x"E2", x"AA", x"64", x"03", x"BC", x"12", x"8C", x"AD", x"9D", x"10", x"16", x"F7", x"00", x"4A", x"AE", x"13", x"35", x"A1", x"43", x"7A", x"83",
  x"74", x"40", x"D9", x"94", x"F8", x"92", x"81", x"45", x"AF", x"C4", x"82", x"45", x"3F", x"37", x"16", x"12", x"A6", x"DB", x"2C", x"03", x"22", x"EA", x"7B", x"F7", x"27",
  x"EF", x"E8", x"A8", x"FE", x"A0", x"A4", x"1D", x"4E", x"31", x"BC", x"A4", x"2E", x"00", x"C4", x"78", x"E5", x"9C", x"D6", x"1F", x"85", x"45", x"6E", x"79", x"AB", x"7C",
  x"A5", x"0A", x"CA", x"6F", x"65", x"F7", x"19", x"D7", x"F0", x"ED", x"8B", x"C0", x"02", x"2F", x"34", x"6B", x"0D", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AB", x"E2", x"AA", x"64", x"03", x"BC", x"12", x"AB", x"94", x"A3",
  x"51", x"28", x"92", x"00", x"41", x"C3", x"BD", x"03", x"31", x"E7", x"B3", x"36", x"7F", x"67", x"2E", x"90", x"DA", x"DD", x"1F", x"EF", x"76", x"A5", x"96", x"8F", x"34",
  x"19", x"30", x"E2", x"AB", x"D3", x"FA", x"B9", x"3E", x"BD", x"49", x"A8", x"4A", x"CE", x"DF", x"69", x"73", x"24", x"41", x"4D", x"1F", x"04", x"B9", x"98", x"C1", x"CA",
  x"5B", x"68", x"3C", x"94", x"C4", x"DC", x"17", x"28", x"1B", x"8E", x"5E", x"78", x"16", x"58", x"1D", x"29", x"EE", x"82", x"67", x"4A", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AB", x"E2", x"AA", x"64", x"03", x"BC", x"12",
  x"15", x"AD", x"4F", x"33", x"EF", x"1F", x"00", x"48", x"1E", x"15", x"89", x"4E", x"FF", x"0A", x"41", x"66", x"E7", x"2F", x"9A", x"F1", x"B0", x"03", x"6B", x"7B", x"71",
  x"19", x"12", x"38", x"DE", x"93", x"96", x"B6", x"08", x"FA", x"4E", x"C7", x"0F", x"42", x"DF", x"BF", x"39", x"0E", x"9F", x"54", x"74", x"F3", x"7A", x"D2", x"A0", x"41",
  x"B6", x"FC", x"E4", x"98", x"5C", x"CB", x"63", x"0E", x"70", x"1D", x"2B", x"DB", x"08", x"66", x"47", x"71", x"43", x"A2", x"43", x"36", x"92", x"DC", x"27", x"B3", x"16",
  x"16", x"4F", x"A7", x"7A", x"D5", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"AA", x"AA", x"AA", x"AA",
  x"AA", x"AA", x"AA", x"AB", x"DC", x"43", x"8E", x"53", x"BA", x"E4", x"62", x"2F", x"1F", x"36", x"F0", x"1D", x"00", x"4D", x"44", x"7F", x"86", x"3A", x"CC", x"18", x"58",
  x"24", x"B3", x"2A", x"79", x"E5", x"6B", x"00", x"F5", x"E5", x"AA", x"BC", x"3D", x"F2", x"35", x"82", x"9F", x"2F", x"80", x"7A", x"19", x"C5", x"2A", x"A0", x"F4", x"0E",
  x"D8", x"E3", x"B1", x"3B", x"4B", x"D9", x"1D", x"83", x"F1", x"09", x"68", x"D1", x"EE", x"C8", x"4F", x"E8", x"75", x"3A", x"BB", x"9C", x"64", x"13", x"F1", x"9C", x"35",
  x"60", x"ED", x"E6", x"B4", x"A1", x"92", x"86", x"3E", x"B3", x"1C", x"BF", x"9E", x"DF", x"FF", x"2A", x"D4", x"B7", x"97", x"66", x"3B", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AB", x"1E", x"C0", x"97", x"39", x"05", x"BD",
  x"15", x"AD", x"4F", x"33", x"EF", x"1F", x"00", x"3D", x"28", x"FA", x"00", x"48", x"9E", x"3E", x"F3", x"53", x"67", x"E0", x"15", x"0D", x"10", x"60", x"9B", x"82", x"76",
  x"DB", x"26", x"CD", x"6B", x"A1", x"5D", x"48", x"12", x"FD", x"57", x"6C", x"F8", x"2E", x"F6", x"C5", x"8E", x"46", x"BA", x"1C", x"1A", x"D3", x"F9", x"1E", x"0D", x"81",
  x"F8", x"2E", x"E9", x"44", x"57", x"E1", x"09", x"1C", x"FC", x"7C", x"AB", x"E8", x"1D", x"D0", x"05", x"6F", x"B9", x"2E", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AB", x"E2", x"AA", x"64", x"03", x"BC", x"12", x"AC",
  x"9D", x"70", x"FA", x"CB", x"F9", x"00", x"4E", x"D0", x"0D", x"CE", x"3A", x"7D", x"33", x"98", x"E2", x"7D", x"8C", x"14", x"7C", x"F5", x"93", x"7E", x"87", x"62", x"06",
  x"35", x"26", x"C3", x"C1", x"F8", x"4A", x"68", x"AC", x"57", x"1F", x"9F", x"E7", x"2F", x"CA", x"A1", x"E6", x"96", x"43", x"27", x"B6", x"86", x"CA", x"5B", x"15", x"C2",
  x"D4", x"9D", x"A2", x"4D", x"F9", x"ED", x"EA", x"9B", x"91", x"3D", x"C8", x"BF", x"10", x"C5", x"DA", x"F6", x"27", x"21", x"A9", x"BE", x"55", x"65", x"D7", x"62", x"FD",
  x"0C", x"08", x"8D", x"F0", x"FE", x"B9", x"1E", x"1C", x"2C", x"0A", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AB", x"E2", x"AA", x"64", x"03", x"BC", x"12", x"B5", x"28", x"56", x"2A", x"FF", x"A3", x"00", x"30", x"73", x"D1",
  x"C2", x"4B", x"F7", x"3E", x"CE", x"11", x"06", x"BB", x"77", x"13", x"02", x"EC", x"74", x"E7", x"37", x"F6", x"64", x"FA", x"0D", x"FF", x"39", x"74", x"84", x"A5", x"A7",
  x"48", x"48", x"A0", x"DF", x"30", x"A0", x"9A", x"7D", x"AF", x"86", x"E0", x"F0", x"0F", x"E0", x"CD", x"B7", x"01", x"7E", x"35", x"AD", x"8D", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AB", x"E2", x"AA", x"64", x"03", x"BC",
  x"12", x"23", x"A3", x"2E", x"1E", x"C5", x"CB", x"00", x"60", x"1C", x"A0", x"3D", x"6F", x"45", x"C1", x"98", x"2A", x"61", x"83", x"FE", x"A6", x"BF", x"55", x"8E", x"0C",
  x"36", x"C2", x"79", x"0A", x"3F", x"42", x"B1", x"42", x"3A", x"26", x"44", x"94", x"E1", x"55", x"51", x"7B", x"FB", x"62", x"1F", x"2C", x"D5", x"D3", x"46", x"C5", x"C7",
  x"64", x"F5", x"65", x"89", x"15", x"26", x"1A", x"64", x"73", x"23", x"0D", x"25", x"6C", x"FE", x"A8", x"EA", x"58", x"73", x"7F", x"E0", x"B9", x"CA", x"A7", x"39", x"9E",
  x"45", x"6B", x"90", x"F5", x"56", x"32", x"78", x"50", x"D6", x"7A", x"43", x"DE", x"1E", x"31", x"41", x"D0", x"7D", x"F1", x"73", x"E5", x"CE", x"D1", x"A2", x"F4", x"1D",
  x"4C", x"4F", x"2B", x"DF", x"17", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"AA", x"AA", x"AA", x"AA",
  x"AA", x"AA", x"AA", x"AB", x"E2", x"AA", x"64", x"03", x"BC", x"12", x"15", x"AD", x"4F", x"33", x"EF", x"1F", x"00", x"4E", x"1A", x"20", x"2C", x"38", x"81", x"F4", x"3A",
  x"96", x"2F", x"7A", x"8B", x"B6", x"89", x"3C", x"1C", x"01", x"86", x"95", x"13", x"DC", x"75", x"1F", x"C5", x"6C", x"54", x"89", x"06", x"CA", x"29", x"FB", x"57", x"15",
  x"DB", x"85", x"8C", x"2A", x"6E", x"29", x"57", x"A5", x"3B", x"B1", x"D5", x"EA", x"02", x"B9", x"2D", x"BD", x"FC", x"63", x"84", x"8A", x"D8", x"33", x"CA", x"D2", x"01",
  x"5F", x"03", x"67", x"49", x"61", x"C2", x"B3", x"BD", x"BB", x"C6", x"01", x"37", x"6B", x"41", x"BC", x"8B", x"13", x"0F", x"E2", x"CD", x"C8", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AB", x"E2", x"AA", x"64", x"03", x"BC",
  x"12", x"15", x"AD", x"4F", x"33", x"EF", x"1F", x"00", x"33", x"D0", x"0C", x"5D", x"31", x"6B", x"B4", x"92", x"B4", x"1B", x"65", x"9E", x"D7", x"3E", x"43", x"68", x"48",
  x"9F", x"4C", x"12", x"04", x"A5", x"E0", x"19", x"9E", x"3C", x"A9", x"56", x"DE", x"EE", x"2D", x"68", x"EE", x"91", x"70", x"61", x"E3", x"D2", x"A1", x"9E", x"85", x"C2",
  x"E4", x"39", x"D7", x"EF", x"71", x"4E", x"B1", x"02", x"CF", x"DF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AB", x"E2", x"AA", x"64", x"03", x"BC", x"12", x"15", x"AD", x"4F", x"33", x"EF", x"1F", x"00", x"4A", x"3B", x"74",
  x"14", x"DE", x"6D", x"82", x"87", x"A3", x"43", x"BB", x"9C", x"2E", x"27", x"3C", x"E7", x"EA", x"65", x"FF", x"15", x"4F", x"A9", x"49", x"2F", x"E3", x"E7", x"E7", x"60",
  x"46", x"96", x"F1", x"04", x"05", x"CE", x"C9", x"A8", x"69", x"40", x"15", x"64", x"87", x"14", x"9D", x"EB", x"E2", x"4E", x"6D", x"A1", x"F7", x"09", x"23", x"1E", x"A1",
  x"69", x"90", x"D9", x"7D", x"43", x"7F", x"0F", x"74", x"69", x"3A", x"24", x"92", x"14", x"18", x"DC", x"1B", x"72", x"91", x"28", x"34", x"07", x"E8", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AB", x"54", x"F6", x"10", x"DD",
  x"AA", x"13", x"54", x"84", x"7B", x"A7", x"12", x"FA", x"00", x"53", x"BE", x"C1", x"E1", x"33", x"AE", x"3E", x"89", x"E4", x"80", x"07", x"67", x"46", x"67", x"1A", x"61",
  x"2B", x"3D", x"14", x"5B", x"F7", x"08", x"0A", x"76", x"BE", x"FB", x"04", x"DB", x"AC", x"54", x"94", x"0C", x"E4", x"45", x"4F", x"AA", x"2F", x"C3", x"A2", x"99", x"B8",
  x"E3", x"4D", x"7C", x"27", x"4F", x"98", x"0A", x"DA", x"EB", x"6E", x"64", x"25", x"0F", x"D9", x"49", x"68", x"AF", x"E7", x"98", x"03", x"C1", x"B3", x"D9", x"50", x"5C",
  x"75", x"55", x"84", x"88", x"E6", x"0B", x"0C", x"DE", x"F5", x"5B", x"3C", x"F4", x"44", x"D0", x"2E", x"B2", x"DB", x"F4", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AB", x"E2", x"AA", x"64", x"03", x"BC", x"12", x"56", x"CD",
  x"FA", x"B4", x"2A", x"EA", x"00", x"5C", x"2B", x"89", x"EF", x"40", x"E0", x"79", x"E1", x"AA", x"C9", x"7F", x"69", x"39", x"9F", x"38", x"2D", x"83", x"19", x"CB", x"6B",
  x"76", x"A0", x"63", x"68", x"F6", x"30", x"4E", x"CB", x"D5", x"88", x"66", x"61", x"83", x"D3", x"F3", x"A0", x"91", x"9F", x"E2", x"1D", x"D5", x"F9", x"41", x"41", x"48",
  x"C8", x"8D", x"75", x"C0", x"B7", x"3F", x"8D", x"DC", x"E4", x"84", x"5B", x"8B", x"A5", x"EE", x"95", x"62", x"69", x"52", x"1B", x"40", x"D2", x"B0", x"2F", x"6A", x"FB",
  x"98", x"67", x"3F", x"14", x"82", x"4F", x"C6", x"01", x"0D", x"C9", x"44", x"69", x"37", x"CC", x"80", x"B6", x"AD", x"64", x"1B", x"22", x"8D", x"58", x"8F", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AB", x"E2", x"AA", x"64",
  x"03", x"BC", x"12", x"15", x"AD", x"4F", x"33", x"EF", x"1F", x"00", x"34", x"09", x"5B", x"D0", x"C3", x"F8", x"8A", x"CC", x"5C", x"BD", x"51", x"8E", x"9C", x"C1", x"D0",
  x"F7", x"1A", x"D1", x"1D", x"59", x"38", x"50", x"B3", x"A8", x"5C", x"B1", x"03", x"E2", x"4E", x"21", x"6A", x"96", x"8A", x"4A", x"85", x"90", x"BD", x"64", x"E8", x"DD",
  x"10", x"3D", x"A9", x"B9", x"E3", x"CB", x"67", x"45", x"C8", x"56", x"86", x"9E", x"A9", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AB", x"23", x"D3", x"EB", x"44", x"69", x"8E", x"15", x"AD", x"4F", x"33", x"EF", x"1F", x"00",
  x"3A", x"61", x"42", x"56", x"A5", x"05", x"42", x"80", x"D4", x"C6", x"CA", x"03", x"61", x"E0", x"18", x"5E", x"C9", x"89", x"97", x"0C", x"93", x"4D", x"C5", x"97", x"62",
  x"D1", x"2E", x"72", x"3F", x"44", x"E3", x"94", x"EE", x"CF", x"C9", x"33", x"3A", x"87", x"04", x"7A", x"92", x"C6", x"BB", x"B9", x"56", x"F7", x"DE", x"F5", x"A4", x"EB",
  x"40", x"2F", x"67", x"5F", x"57", x"91", x"73", x"FD", x"23", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AB", x"E2", x"AA", x"64", x"03", x"BC", x"12", x"AE", x"EE", x"64", x"5F", x"DF", x"D0", x"00", x"5B", x"8A", x"1E", x"2B",
  x"7F", x"5D", x"6E", x"F0", x"25", x"47", x"DC", x"DE", x"75", x"5C", x"40", x"AA", x"12", x"F6", x"2B", x"B8", x"DC", x"9E", x"AB", x"47", x"9E", x"77", x"84", x"CC", x"01",
  x"BA", x"16", x"AA", x"03", x"10", x"4A", x"9F", x"46", x"4D", x"3C", x"33", x"8E", x"AC", x"C2", x"13", x"A6", x"7C", x"A0", x"A9", x"46", x"5E", x"10", x"06", x"C8", x"D4",
  x"3E", x"6C", x"20", x"C0", x"3E", x"32", x"88", x"E9", x"8F", x"D9", x"14", x"3C", x"46", x"7F", x"10", x"F6", x"5E", x"10", x"D2", x"F1", x"48", x"12", x"27", x"20", x"4E",
  x"C4", x"CD", x"D0", x"76", x"F6", x"DB", x"F0", x"29", x"65", x"C5", x"1B", x"9C", x"86", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AB", x"E2", x"AA", x"64", x"03", x"BC", x"12", x"62", x"C9", x"54", x"C0", x"43", x"CB", x"00",
  x"2E", x"2A", x"39", x"C0", x"7F", x"BE", x"9D", x"81", x"A3", x"37", x"D5", x"0B", x"80", x"F6", x"BD", x"53", x"6E", x"1C", x"D8", x"B7", x"E8", x"D9", x"3D", x"CD", x"30",
  x"B0", x"11", x"BC", x"62", x"DD", x"48", x"4F", x"4C", x"0B", x"53", x"B1", x"0A", x"FA", x"0F", x"89", x"76", x"EE", x"78", x"68", x"23", x"A9", x"D3", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AB", x"E2", x"AA", x"64", x"03",
  x"BC", x"12", x"E1", x"B8", x"D8", x"31", x"A5", x"BC", x"00", x"59", x"44", x"52", x"04", x"0F", x"79", x"79", x"6E", x"12", x"4E", x"28", x"A7", x"76", x"6D", x"84", x"11",
  x"07", x"29", x"17", x"71", x"55", x"9C", x"63", x"44", x"E1", x"60", x"59", x"14", x"78", x"CB", x"F5", x"09", x"94", x"90", x"D2", x"B6", x"C9", x"3B", x"0D", x"51", x"13",
  x"34", x"B0", x"6C", x"4C", x"C3", x"AC", x"A4", x"2F", x"BA", x"3C", x"EA", x"A8", x"C1", x"12", x"FD", x"33", x"43", x"AB", x"05", x"EF", x"E2", x"2A", x"1E", x"2C", x"3B",
  x"26", x"61", x"E9", x"B5", x"03", x"2D", x"6A", x"FD", x"4E", x"85", x"CD", x"75", x"C3", x"11", x"DF", x"33", x"31", x"03", x"16", x"51", x"74", x"A8", x"F2", x"5F", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AB", x"E2", x"AA",
  x"64", x"03", x"BC", x"12", x"1E", x"22", x"3D", x"C4", x"76", x"5C", x"00", x"35", x"6E", x"01", x"76", x"7D", x"05", x"3C", x"18", x"56", x"7F", x"CA", x"C7", x"00", x"2D",
  x"6F", x"DF", x"DB", x"D7", x"6E", x"DA", x"E9", x"92", x"EB", x"8C", x"4A", x"27", x"7A", x"D1", x"FD", x"88", x"D3", x"FA", x"A0", x"28", x"02", x"EA", x"81", x"10", x"03",
  x"36", x"03", x"B4", x"07", x"21", x"B2", x"86", x"0B", x"58", x"17", x"D9", x"DF", x"D7", x"EC", x"44", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AB", x"E2", x"AA", x"64", x"03", x"BC", x"12", x"15", x"AD", x"4F", x"33", x"EF",
  x"1F", x"00", x"60", x"95", x"CD", x"46", x"8C", x"E4", x"76", x"F5", x"65", x"A9", x"01", x"AB", x"BA", x"33", x"F3", x"63", x"A1", x"D8", x"7D", x"B6", x"B2", x"20", x"9B",
  x"E5", x"26", x"5A", x"5F", x"6D", x"2A", x"DF", x"C9", x"65", x"AC", x"B2", x"AA", x"78", x"3F", x"5F", x"0D", x"19", x"38", x"BF", x"EE", x"A1", x"4F", x"2E", x"C0", x"4A",
  x"68", x"9B", x"41", x"CD", x"3D", x"E8", x"F1", x"1F", x"15", x"1D", x"37", x"AB", x"0C", x"27", x"7C", x"86", x"A5", x"B1", x"24", x"4D", x"FA", x"D9", x"E2", x"47", x"92",
  x"9B", x"9E", x"8A", x"6F", x"4A", x"4E", x"63", x"23", x"FA", x"FF", x"4B", x"44", x"6E", x"FF", x"F7", x"91", x"D1", x"83", x"DC", x"51", x"E9", x"EF", x"3A", x"0C", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AB", x"94", x"ED",
  x"52", x"E7", x"46", x"CF", x"07", x"D4", x"E9", x"01", x"02", x"4C", x"00", x"4F", x"41", x"6F", x"CE", x"D2", x"84", x"06", x"03", x"7F", x"0A", x"45", x"0A", x"83", x"CC",
  x"BD", x"DF", x"77", x"A5", x"74", x"B9", x"9E", x"94", x"87", x"23", x"95", x"D4", x"74", x"94", x"9E", x"27", x"47", x"89", x"40", x"8F", x"B7", x"08", x"E9", x"8D", x"BB",
  x"19", x"08", x"17", x"1D", x"6A", x"32", x"AD", x"13", x"BD", x"07", x"FC", x"74", x"A5", x"CF", x"3F", x"C9", x"55", x"4C", x"DA", x"A8", x"DC", x"92", x"C7", x"5F", x"E1",
  x"6C", x"5D", x"61", x"8E", x"3A", x"C9", x"00", x"5A", x"9E", x"DC", x"38", x"E9", x"11", x"47", x"12", x"0E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AB", x"EA", x"05", x"0B", x"55", x"25", x"33", x"15", x"AD", x"4F", x"33",
  x"EF", x"1F", x"00", x"4A", x"9C", x"DE", x"FF", x"2B", x"00", x"81", x"02", x"AA", x"42", x"E7", x"9C", x"0D", x"AA", x"D5", x"01", x"CA", x"7A", x"AD", x"C3", x"11", x"16",
  x"D4", x"47", x"E6", x"36", x"E6", x"FF", x"2E", x"4F", x"10", x"CE", x"34", x"56", x"87", x"38", x"56", x"CD", x"91", x"0E", x"0F", x"13", x"0A", x"34", x"A9", x"18", x"66",
  x"34", x"01", x"14", x"5D", x"EC", x"26", x"5D", x"6D", x"FA", x"FD", x"B1", x"52", x"0B", x"A7", x"E4", x"B4", x"E6", x"D9", x"DD", x"C6", x"4A", x"11", x"74", x"08", x"E7",
  x"77", x"93", x"5E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA",
  x"AA", x"AB", x"E2", x"AA", x"64", x"03", x"BC", x"12", x"15", x"AD", x"4F", x"33", x"EF", x"1F", x"00", x"5B", x"58", x"F3", x"98", x"B0", x"13", x"A3", x"52", x"24", x"62",
  x"F7", x"6F", x"24", x"14", x"64", x"02", x"87", x"1B", x"3E", x"13", x"19", x"54", x"0C", x"01", x"AB", x"BE", x"FB", x"2A", x"60", x"67", x"11", x"67", x"F5", x"A7", x"DD",
  x"14", x"99", x"46", x"18", x"10", x"08", x"7F", x"0C", x"03", x"46", x"04", x"E0", x"63", x"C9", x"3E", x"AA", x"64", x"90", x"56", x"64", x"5D", x"4E", x"7E", x"26", x"8F",
  x"BF", x"4A", x"CC", x"37", x"48", x"62", x"04", x"9A", x"71", x"AD", x"6E", x"3E", x"91", x"68", x"7F", x"EB", x"CB", x"E4", x"72", x"6C", x"68", x"F7", x"BF", x"88", x"0E",
  x"00", x"3E", x"0C", x"B0", x"BB", x"DA", x"57", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"AA", x"AA",
  x"AA", x"AA", x"AA", x"AA", x"AA", x"AB", x"E2", x"AA", x"64", x"03", x"BC", x"12", x"0F", x"ED", x"B0", x"37", x"02", x"3A", x"00", x"58", x"4A", x"82", x"20", x"B4", x"FD",
  x"B8", x"1A", x"02", x"0D", x"6E", x"12", x"5E", x"8B", x"63", x"F1", x"22", x"EB", x"0B", x"75", x"1E", x"2E", x"A0", x"A7", x"D5", x"AF", x"63", x"65", x"BD", x"06", x"E9",
  x"13", x"DF", x"DF", x"BF", x"88", x"52", x"3D", x"BE", x"DE", x"91", x"89", x"1E", x"98", x"74", x"2E", x"AC", x"68", x"71", x"CA", x"35", x"B5", x"1F", x"FA", x"71", x"01",
  x"9D", x"BD", x"C0", x"FE", x"C0", x"AB", x"B6", x"4C", x"9A", x"F9", x"AF", x"02", x"C3", x"65", x"A9", x"39", x"B6", x"49", x"9D", x"DB", x"C3", x"0E", x"29", x"9D", x"E4",
  x"CA", x"AC", x"FB", x"EC", x"9E", x"6E", x"4E", x"6E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"AA",
  x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AB", x"66", x"20", x"B6", x"80", x"AF", x"AD", x"D6", x"75", x"38", x"6F", x"24", x"9A", x"00", x"52", x"96", x"D0", x"CE", x"60",
  x"32", x"CE", x"C7", x"19", x"E9", x"7D", x"4B", x"6E", x"B2", x"8D", x"27", x"D8", x"A7", x"97", x"99", x"DE", x"E4", x"2A", x"B7", x"5C", x"4E", x"AA", x"E0", x"B7", x"8E",
  x"B7", x"88", x"29", x"23", x"B9", x"FB", x"92", x"D6", x"96", x"EE", x"13", x"8A", x"5B", x"36", x"D2", x"58", x"76", x"FE", x"15", x"C8", x"30", x"61", x"58", x"CF", x"4E",
  x"0B", x"DF", x"68", x"CB", x"78", x"BF", x"DF", x"0A", x"F0", x"45", x"B8", x"8D", x"53", x"86", x"B0", x"DF", x"E1", x"E2", x"BB", x"52", x"73", x"72", x"A1", x"A3", x"96",
  x"D7", x"66", x"B8", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA",
  x"AA", x"AB", x"E2", x"AA", x"64", x"03", x"BC", x"12", x"4A", x"0E", x"C0", x"EE", x"14", x"44", x"00", x"5A", x"A3", x"F2", x"79", x"50", x"9A", x"F6", x"13", x"4C", x"6B",
  x"40", x"8E", x"09", x"07", x"DF", x"56", x"31", x"17", x"10", x"0F", x"22", x"5D", x"6E", x"98", x"2C", x"96", x"78", x"90", x"B5", x"31", x"9E", x"C1", x"32", x"ED", x"4B",
  x"1F", x"1F", x"A4", x"CD", x"B6", x"E5", x"28", x"12", x"20", x"E7", x"90", x"84", x"E5", x"95", x"83", x"A1", x"04", x"96", x"DF", x"6A", x"5F", x"8B", x"BE", x"7D", x"63",
  x"69", x"B2", x"0E", x"8B", x"03", x"AA", x"8B", x"0C", x"C4", x"F9", x"BF", x"F5", x"3D", x"97", x"CE", x"F7", x"CD", x"13", x"A2", x"18", x"DD", x"B5", x"35", x"34", x"C1",
  x"E0", x"AD", x"71", x"EA", x"48", x"B2", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"AA", x"AA", x"AA",
  x"AA", x"AA", x"AA", x"AA", x"AB", x"F8", x"54", x"66", x"88", x"02", x"3C", x"15", x"AD", x"4F", x"33", x"EF", x"1F", x"00", x"40", x"4B", x"D1", x"E4", x"B0", x"EB", x"B0",
  x"37", x"31", x"18", x"D9", x"54", x"FC", x"28", x"30", x"04", x"CD", x"F7", x"CF", x"3E", x"D9", x"DF", x"43", x"98", x"95", x"20", x"64", x"2E", x"B3", x"C7", x"65", x"4C",
  x"F9", x"01", x"A6", x"63", x"EA", x"86", x"20", x"4C", x"46", x"64", x"9E", x"E7", x"D2", x"8F", x"76", x"AB", x"31", x"26", x"80", x"7E", x"FB", x"4F", x"E4", x"D4", x"F3",
  x"B8", x"0A", x"D1", x"02", x"62", x"2A", x"58", x"81", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"AA",
  x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AB", x"E2", x"AA", x"64", x"03", x"BC", x"12", x"FA", x"30", x"53", x"4A", x"B0", x"C2", x"00", x"63", x"88", x"25", x"0F", x"1A",
  x"83", x"FC", x"A6", x"3C", x"DB", x"10", x"37", x"89", x"C3", x"28", x"44", x"A9", x"D8", x"D5", x"95", x"C8", x"C6", x"63", x"03", x"A8", x"B9", x"BC", x"30", x"A6", x"E4",
  x"36", x"37", x"B2", x"63", x"6B", x"10", x"B4", x"49", x"34", x"12", x"2C", x"F3", x"19", x"9A", x"88", x"5C", x"03", x"54", x"DE", x"AC", x"4E", x"2E", x"96", x"BB", x"65",
  x"3B", x"59", x"6C", x"10", x"A8", x"F4", x"92", x"25", x"0B", x"EB", x"55", x"75", x"2A", x"B9", x"27", x"15", x"EA", x"D4", x"5A", x"DA", x"A8", x"FB", x"79", x"8B", x"9F",
  x"40", x"AA", x"60", x"7F", x"1F", x"8C", x"FE", x"94", x"F4", x"4E", x"E5", x"E6", x"A0", x"95", x"0F", x"04", x"21", x"2B", x"DD", x"45", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AB", x"E2", x"AA", x"64", x"03", x"BC", x"12",
  x"16", x"A6", x"88", x"7A", x"34", x"DA", x"00", x"3D", x"F5", x"4B", x"97", x"09", x"77", x"96", x"D5", x"9B", x"C3", x"15", x"5A", x"FE", x"1D", x"33", x"C2", x"91", x"7B",
  x"9A", x"2A", x"2F", x"DB", x"46", x"D8", x"B5", x"C1", x"08", x"0C", x"73", x"CA", x"07", x"74", x"66", x"10", x"CE", x"55", x"B6", x"1B", x"74", x"1A", x"B7", x"44", x"45",
  x"6C", x"04", x"42", x"CF", x"E2", x"17", x"32", x"C7", x"3F", x"61", x"13", x"5B", x"07", x"D7", x"89", x"0B", x"8F", x"BB", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AB", x"69", x"10", x"9B", x"F5", x"08", x"BA", x"15",
  x"AD", x"4F", x"33", x"EF", x"1F", x"00", x"4B", x"F4", x"74", x"D7", x"EC", x"6E", x"20", x"22", x"79", x"94", x"D4", x"35", x"E7", x"04", x"46", x"4A", x"37", x"37", x"3F",
  x"08", x"6A", x"69", x"07", x"05", x"6D", x"77", x"03", x"12", x"9C", x"0A", x"D9", x"20", x"A1", x"B0", x"D6", x"A1", x"31", x"6A", x"24", x"E3", x"94", x"EA", x"57", x"19",
  x"F6", x"50", x"5F", x"DB", x"D1", x"89", x"F7", x"38", x"84", x"D3", x"CF", x"82", x"6B", x"B3", x"22", x"B4", x"17", x"02", x"AB", x"73", x"59", x"18", x"23", x"20", x"44",
  x"93", x"13", x"67", x"FD", x"76", x"BD", x"70", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"AA", x"AA",
  x"AA", x"AA", x"AA", x"AA", x"AA", x"AB", x"E2", x"AA", x"64", x"03", x"BC", x"12", x"15", x"AD", x"4F", x"33", x"EF", x"1F", x"00", x"62", x"FD", x"8D", x"C6", x"8A", x"CA",
  x"04", x"7D", x"84", x"0C", x"39", x"9C", x"A7", x"91", x"15", x"9F", x"F7", x"95", x"E9", x"72", x"0A", x"B3", x"EF", x"6D", x"C3", x"BD", x"39", x"E3", x"4B", x"BA", x"B7",
  x"3E", x"FF", x"FD", x"32", x"8F", x"FA", x"09", x"B0", x"9A", x"C5", x"73", x"10", x"55", x"D8", x"09", x"3F", x"38", x"B1", x"2D", x"5C", x"0B", x"09", x"E9", x"E6", x"54",
  x"8F", x"79", x"83", x"84", x"C7", x"D0", x"22", x"5D", x"5F", x"44", x"63", x"31", x"E6", x"4E", x"0A", x"14", x"96", x"93", x"F7", x"C9", x"DF", x"3D", x"E2", x"14", x"CE",
  x"8D", x"32", x"36", x"48", x"DB", x"FF", x"78", x"D5", x"9A", x"1B", x"E3", x"F5", x"10", x"38", x"A9", x"03", x"8E", x"D7", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AB", x"E1", x"59", x"F5", x"46", x"2F", x"98", x"15", x"AD",
  x"4F", x"33", x"EF", x"1F", x"00", x"3E", x"81", x"96", x"F3", x"02", x"B0", x"B4", x"FB", x"00", x"A3", x"D2", x"50", x"6E", x"31", x"45", x"2C", x"15", x"10", x"94", x"3E",
  x"94", x"96", x"77", x"F6", x"0A", x"BF", x"51", x"C5", x"89", x"D9", x"8A", x"FB", x"2D", x"F4", x"48", x"DC", x"2E", x"42", x"29", x"5A", x"90", x"FC", x"F9", x"B5", x"E9",
  x"1C", x"AE", x"D3", x"39", x"E2", x"B3", x"9A", x"65", x"64", x"5B", x"85", x"62", x"D0", x"8F", x"E2", x"00", x"C7", x"FD", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AB", x"7E", x"8F", x"13", x"B1", x"B6", x"1E", x"15", x"AD",
  x"4F", x"33", x"EF", x"1F", x"00", x"44", x"C5", x"2D", x"15", x"EF", x"95", x"BB", x"AC", x"33", x"93", x"49", x"29", x"1E", x"B3", x"00", x"F0", x"D7", x"0F", x"3A", x"8B",
  x"CB", x"8D", x"A5", x"10", x"4D", x"A1", x"64", x"AF", x"B9", x"19", x"E3", x"C2", x"CA", x"81", x"34", x"D6", x"E2", x"A4", x"CB", x"7F", x"84", x"5C", x"38", x"92", x"B2",
  x"6B", x"F9", x"EF", x"3F", x"99", x"B7", x"D4", x"01", x"3E", x"9B", x"5F", x"0D", x"76", x"30", x"63", x"7B", x"C6", x"E2", x"A0", x"DF", x"3B", x"CA", x"78", x"13", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AB", x"E2", x"AA",
  x"64", x"03", x"BC", x"12", x"8B", x"AB", x"AD", x"37", x"3F", x"E4", x"00", x"52", x"BE", x"0B", x"DD", x"CD", x"5A", x"59", x"B5", x"47", x"6B", x"C5", x"49", x"42", x"D9",
  x"12", x"83", x"F6", x"5A", x"B2", x"AA", x"8E", x"E4", x"92", x"A6", x"FD", x"E1", x"6E", x"40", x"E4", x"E0", x"FD", x"C5", x"B8", x"C0", x"9E", x"E1", x"68", x"94", x"7A",
  x"E9", x"44", x"B1", x"E0", x"6C", x"37", x"44", x"19", x"21", x"65", x"32", x"5B", x"7A", x"D1", x"D4", x"7F", x"2D", x"BB", x"71", x"4F", x"27", x"9B", x"A3", x"C7", x"84",
  x"23", x"56", x"C4", x"09", x"EB", x"3C", x"24", x"7C", x"52", x"F0", x"D9", x"7A", x"93", x"79", x"EF", x"A6", x"72", x"B0", x"CD", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AB", x"E2", x"AA", x"64", x"03", x"BC", x"12", x"15",
  x"AD", x"4F", x"33", x"EF", x"1F", x"00", x"3C", x"90", x"11", x"F4", x"71", x"A5", x"EB", x"9D", x"44", x"11", x"90", x"D0", x"A5", x"D5", x"0A", x"18", x"FE", x"CD", x"62",
  x"52", x"0C", x"4C", x"DB", x"87", x"05", x"3F", x"BF", x"01", x"F1", x"96", x"2D", x"BA", x"EF", x"C3", x"4D", x"D8", x"D1", x"77", x"FD", x"09", x"90", x"AE", x"8A", x"F5",
  x"64", x"EE", x"29", x"EF", x"B8", x"B7", x"61", x"B0", x"3E", x"BC", x"91", x"45", x"DE", x"37", x"8E", x"3C", x"EE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AB", x"4D", x"3A", x"F6", x"79", x"60", x"AF", x"1D", x"DD", x"9F",
  x"ED", x"CD", x"33", x"00", x"43", x"20", x"0D", x"65", x"5B", x"78", x"B4", x"E2", x"44", x"30", x"48", x"95", x"0A", x"AB", x"85", x"E1", x"96", x"8F", x"E4", x"59", x"E8",
  x"6A", x"7C", x"7E", x"34", x"F3", x"6E", x"52", x"E1", x"DB", x"D2", x"B2", x"85", x"F0", x"FB", x"4E", x"00", x"CC", x"B8", x"E4", x"A7", x"33", x"17", x"9C", x"00", x"C0",
  x"30", x"AA", x"46", x"0B", x"6B", x"D2", x"EB", x"54", x"1C", x"BF", x"D9", x"60", x"3B", x"7B", x"69", x"DA", x"44", x"24", x"02", x"AB", x"E5", x"8C", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AB", x"E2", x"AA", x"64", x"03",
  x"BC", x"12", x"15", x"AD", x"4F", x"33", x"EF", x"1F", x"00", x"3A", x"CC", x"5C", x"42", x"AF", x"CC", x"07", x"AD", x"20", x"7E", x"BA", x"68", x"30", x"D4", x"06", x"A7",
  x"CD", x"13", x"27", x"01", x"F3", x"F5", x"93", x"64", x"22", x"2F", x"9F", x"E8", x"11", x"9B", x"7F", x"0D", x"F4", x"4A", x"3C", x"7D", x"E2", x"EE", x"98", x"7A", x"AC",
  x"54", x"3D", x"BD", x"1D", x"B2", x"BA", x"56", x"77", x"CA", x"DA", x"06", x"FC", x"21", x"38", x"F8", x"3A", x"E6", x"8F", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AB", x"E2", x"AA", x"64", x"03", x"BC", x"12", x"15", x"AD",
  x"4F", x"33", x"EF", x"1F", x"00", x"48", x"A1", x"02", x"97", x"2E", x"BE", x"4F", x"BA", x"D1", x"D9", x"71", x"80", x"26", x"20", x"38", x"4C", x"30", x"F4", x"EC", x"42",
  x"C2", x"BE", x"0A", x"F6", x"7F", x"E9", x"2C", x"D8", x"F2", x"AF", x"70", x"A5", x"8F", x"F5", x"F6", x"4E", x"37", x"12", x"F8", x"19", x"42", x"6F", x"23", x"88", x"62",
  x"60", x"49", x"8D", x"82", x"08", x"02", x"B5", x"78", x"34", x"ED", x"9A", x"E8", x"9D", x"90", x"81", x"47", x"9A", x"BD", x"BE", x"5F", x"4A", x"87", x"56", x"97", x"FE",
  x"E0", x"8F", x"4F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA",
  x"AA", x"AB", x"E2", x"AA", x"64", x"03", x"BC", x"12", x"15", x"AD", x"4F", x"33", x"EF", x"1F", x"00", x"50", x"F0", x"C7", x"E5", x"02", x"F3", x"06", x"B3", x"E5", x"D9",
  x"B2", x"70", x"97", x"ED", x"B1", x"7A", x"89", x"61", x"25", x"B3", x"64", x"EB", x"4A", x"1E", x"9A", x"CD", x"26", x"2C", x"49", x"24", x"7A", x"12", x"2B", x"F3", x"80",
  x"66", x"51", x"B7", x"5E", x"86", x"D9", x"5F", x"35", x"AA", x"95", x"EB", x"12", x"AC", x"33", x"15", x"57", x"BE", x"D0", x"64", x"D8", x"A3", x"5C", x"A5", x"60", x"E0",
  x"6D", x"F2", x"A5", x"9F", x"9F", x"FF", x"AA", x"CA", x"A6", x"68", x"FF", x"EA", x"C1", x"40", x"F7", x"47", x"F4", x"F9", x"B6", x"BA", x"58", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AB", x"72", x"19", x"D9", x"9F", x"7E",
  x"B3", x"15", x"AD", x"4F", x"33", x"EF", x"1F", x"00", x"4C", x"1F", x"AF", x"B3", x"EA", x"D8", x"CC", x"A6", x"3F", x"F7", x"07", x"39", x"9E", x"2F", x"FE", x"80", x"E2",
  x"EC", x"93", x"16", x"13", x"46", x"C5", x"A4", x"86", x"4A", x"02", x"99", x"03", x"97", x"ED", x"78", x"62", x"F8", x"A7", x"AD", x"9A", x"3E", x"F4", x"79", x"95", x"53",
  x"F2", x"CC", x"62", x"48", x"8B", x"3B", x"6D", x"92", x"FE", x"97", x"55", x"A6", x"07", x"E7", x"CD", x"85", x"7B", x"5A", x"16", x"58", x"B1", x"EE", x"5F", x"B6", x"37",
  x"38", x"D5", x"62", x"22", x"4E", x"43", x"5D", x"98", x"01", x"5D", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AB", x"E2", x"AA", x"64", x"03", x"BC", x"12", x"5A", x"A9", x"69", x"BC", x"E4", x"DC", x"00", x"30", x"A3", x"89",
  x"3F", x"04", x"93", x"3C", x"AA", x"21", x"92", x"39", x"AC", x"63", x"7F", x"73", x"EC", x"AB", x"B9", x"5D", x"CC", x"8B", x"89", x"99", x"B9", x"2C", x"8C", x"4B", x"A8",
  x"77", x"39", x"B0", x"AB", x"D2", x"DD", x"29", x"67", x"52", x"75", x"D3", x"C7", x"E4", x"86", x"FE", x"DA", x"D1", x"47", x"4E", x"86", x"61", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AB", x"E2", x"AA", x"64", x"03", x"BC",
  x"12", x"15", x"AD", x"4F", x"33", x"EF", x"1F", x"00", x"41", x"71", x"D8", x"6F", x"AE", x"44", x"41", x"E8", x"6A", x"40", x"23", x"5B", x"26", x"71", x"C9", x"59", x"65",
  x"CE", x"2A", x"89", x"EB", x"E9", x"7F", x"9A", x"A7", x"E2", x"06", x"6D", x"DC", x"95", x"C6", x"4A", x"EB", x"2E", x"44", x"3C", x"3D", x"BC", x"E4", x"96", x"76", x"48",
  x"C8", x"C4", x"6B", x"B4", x"8E", x"CA", x"D1", x"58", x"BF", x"8D", x"9E", x"60", x"8D", x"EE", x"B6", x"6D", x"7A", x"4C", x"22", x"99", x"30", x"97", x"08", x"AA", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AB", x"E2", x"AA",
  x"64", x"03", x"BC", x"12", x"2D", x"76", x"B9", x"74", x"28", x"52", x"00", x"62", x"CC", x"23", x"F8", x"CC", x"A2", x"E2", x"E8", x"66", x"20", x"51", x"C6", x"03", x"A0",
  x"7F", x"CE", x"54", x"4C", x"E3", x"0F", x"66", x"80", x"B6", x"E2", x"5D", x"3B", x"A1", x"DD", x"DE", x"B3", x"8B", x"23", x"78", x"CF", x"DB", x"B5", x"22", x"E5", x"E1",
  x"3D", x"C4", x"B9", x"E2", x"14", x"CA", x"02", x"06", x"C0", x"E5", x"1A", x"FF", x"60", x"7E", x"34", x"D2", x"8F", x"49", x"A7", x"5D", x"8D", x"C5", x"0A", x"98", x"64",
  x"CA", x"77", x"FD", x"02", x"67", x"6A", x"4B", x"98", x"44", x"96", x"88", x"51", x"44", x"A7", x"EB", x"6E", x"46", x"0B", x"6C", x"59", x"55", x"8B", x"13", x"E0", x"D2",
  x"AF", x"08", x"11", x"1D", x"09", x"52", x"86", x"6D", x"AE", x"97", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AB", x"B0", x"2E", x"23", x"3E", x"FE", x"00", x"15", x"AD", x"4F", x"33", x"EF", x"1F", x"00", x"5C", x"06", x"53",
  x"D5", x"4D", x"EE", x"7D", x"20", x"27", x"B7", x"BF", x"65", x"8D", x"1F", x"70", x"A8", x"49", x"DD", x"B4", x"70", x"C1", x"CE", x"47", x"F3", x"2C", x"BD", x"28", x"88",
  x"F5", x"39", x"D6", x"30", x"61", x"32", x"E6", x"42", x"C4", x"FC", x"F9", x"E5", x"35", x"E3", x"AA", x"47", x"F6", x"71", x"B0", x"30", x"CF", x"03", x"D2", x"2E", x"05",
  x"BD", x"AB", x"54", x"45", x"FE", x"30", x"1C", x"8E", x"B4", x"1D", x"0E", x"5B", x"11", x"A0", x"B2", x"70", x"9F", x"F0", x"83", x"C9", x"E7", x"8E", x"36", x"AE", x"97",
  x"51", x"E2", x"9F", x"20", x"59", x"41", x"EB", x"5C", x"FB", x"77", x"14", x"7D", x"80", x"FF", x"02", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AB", x"E2", x"AA", x"64", x"03", x"BC", x"12", x"15", x"AD", x"4F", x"33", x"EF",
  x"1F", x"00", x"5A", x"99", x"5D", x"DB", x"04", x"D4", x"A3", x"30", x"27", x"AB", x"3B", x"D7", x"77", x"48", x"F3", x"9C", x"21", x"46", x"E8", x"59", x"CF", x"2F", x"95",
  x"D2", x"6F", x"12", x"CC", x"87", x"12", x"15", x"D3", x"6A", x"C9", x"12", x"56", x"16", x"59", x"56", x"AA", x"88", x"6A", x"1E", x"CE", x"C6", x"63", x"8A", x"8D", x"82",
  x"3D", x"EF", x"E4", x"B2", x"57", x"50", x"2B", x"90", x"90", x"7E", x"10", x"C3", x"22", x"48", x"DF", x"AF", x"33", x"F4", x"C3", x"FE", x"A7", x"B6", x"97", x"B7", x"6D",
  x"13", x"85", x"6C", x"D8", x"01", x"7A", x"6C", x"4F", x"4A", x"A1", x"ED", x"1E", x"CA", x"72", x"B7", x"8C", x"C5", x"B7", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"AB", x"E2", x"AA", x"64", x"03", x"BC", x"12", x"F6", x"E5",
  x"CE", x"75", x"61", x"B7", x"00", x"4B", x"83", x"A2", x"40", x"D7", x"28", x"E5", x"48", x"8E", x"B2", x"CE", x"0A", x"FE", x"B0", x"5C", x"79", x"E1", x"ED", x"3C", x"77",
  x"0F", x"E1", x"9F", x"74", x"3B", x"E0", x"24", x"16", x"73", x"F7", x"C4", x"88", x"7A", x"A8", x"E8", x"7D", x"29", x"C4", x"64", x"68", x"BF", x"E8", x"4F", x"F4", x"18",
  x"DA", x"C8", x"18", x"76", x"BE", x"78", x"F1", x"CD", x"AB", x"08", x"78", x"65", x"02", x"60", x"DC", x"A6", x"B0", x"E6", x"33", x"C5", x"CC", x"8C", x"66", x"05", x"77",
  x"4B", x"1E", x"AB", x"66", x"33", x"33", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
  x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00");
end package;
 
package body util_pkg is
 
	function log2c(n : integer) return integer is
		variable m, p : integer;
	begin
		m := 0;
		p := 1;
		while p < n loop
			m := m + 1;
			p := p * 2;
		end loop;
		return m;
	end function;

end package body;
